LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY FREQDIVN IS
  PORT (
    CLK : IN STD_LOGIC;
    CLK10, CLK100 : OUT STD_LOGIC);
END FREQDIVN;
ARCHITECTURE BEHAVE OF FREQDIVN IS
	SIGNAL X : STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL Y : STD_LOGIC_VECTOR(6 DOWNTO 0);
BEGIN
	PROCESS (CLK)
	BEGIN
		IF (CLK = '1' AND CLK'EVENT) THEN
			IF (X = "1001") THEN
				X <= "0000";
				CLK10 <= '1';
			ELSE
				X <= X + '1';
				CLK10 <= '0';
			END IF;
			IF (Y = "1100100") THEN
				Y <= "0000000";
				CLK100 <= '1';
			ELSE
				Y <= Y + '1';
				CLK100 <= '0';
			END IF;
		END IF;
	END PROCESS;
END BEHAVE;