LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY MYCLOCK IS
	PORT (
		CLK : IN STD_LOGIC;
		EN : IN STD_LOGIC;
		CLR : IN STD_LOGIC;
		VOCOUT : OUT STD_LOGIC;
		SELOUT : OUT STD_LOGIC_VECTOR (0 TO 7);
		DISOUT : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
	);
END MYCLOCK;
ARCHITECTURE BEHAVE OF MYCLOCK IS
	SIGNAL SECONDCO : STD_LOGIC;
	SIGNAL MINUTECO : STD_LOGIC;
	SIGNAL SEL : STD_LOGIC_VECTOR (2 DOWNTO 0);
	SIGNAL DISMUX : STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL CLK_10 : STD_LOGIC;
	SIGNAL CLK_100 : STD_LOGIC;
	SIGNAL SE1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL SE0 : STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL MI1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL MI0 : STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL HO1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL HO0 : STD_LOGIC_VECTOR (3 DOWNTO 0);
	COMPONENT STATECYCLE
		PORT (
			CLK : IN STD_LOGIC;
			CYCOUT : OUT STD_LOGIC_VECTOR(2 DOWNTO 0));
	END COMPONENT;
	COMPONENT DECODE138
		PORT (
			DIN : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
			DOUT : OUT STD_LOGIC_VECTOR (0 TO 7));
	END COMPONENT;
	COMPONENT DISPLAYDECOD
		PORT (
			NUM : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			DISPLAYOUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
	END COMPONENT;

	COMPONENT SECOND
		PORT (
			CLK, EN, CLR : IN STD_LOGIC;
			SEC1, SEC0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			CO : OUT STD_LOGIC);
	END COMPONENT;
	COMPONENT MINUTE
		PORT (
			CLK, EN, CLR : IN STD_LOGIC;
			MIN1, MIN0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			CO : OUT STD_LOGIC);
	END COMPONENT;
	COMPONENT HOUR
		PORT (
			CLK, EN, CLR : IN STD_LOGIC;
			HOU1, HOU0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
	END COMPONENT;
	COMPONENT MUX6
		PORT (
			NUM0, NUM1, NUM2, NUM3, NUM4, NUM5 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			SEL : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			MUX6OUT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
	END COMPONENT;
	COMPONENT FREQDIVN
		PORT (
			CLK : IN STD_LOGIC;
			CLK10, CLK100 : OUT STD_LOGIC);
	END COMPONENT;
	COMPONENT TIMEKEEP
		PORT (
			CLK, CLK1 : IN STD_LOGIC;
			M0, M1, S0, S1 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			TIMEOUT : OUT STD_LOGIC);
	END COMPONENT;
BEGIN
	U1 : TIMEKEEP PORT MAP(CLK, CLK_10, MI1, MI0, SE1, SE0, VOCOUT);
	U2 : FREQDIVN PORT MAP(CLK, CLK_10, CLK_100);
	U3 : SECOND PORT MAP(CLK_100, EN, CLR, SE1, SE0, SECONDCO);
	U4 : MINUTE PORT MAP(SECONDCO, EN, CLR, MI1, MI0, MINUTECO);
	U5 : HOUR PORT MAP(MINUTECO, EN, CLR, HO1, HO0);
	U6 : STATECYCLE PORT MAP(CLK_100, SEL);
	U7 : DECODE138 PORT MAP(SEL, SELOUT);
	U8 : DISPLAYDECOD PORT MAP(DISMUX, DISOUT);
	U9 : MUX6 PORT MAP(HO1, HO0, MI1, MI0, SE1, SE0, SEL, DISMUX);
END BEHAVE;