LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY MINUTE IS
	PORT (
		CLK, EN, CLR : IN STD_LOGIC;
		MIN1, MIN0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		CO : OUT STD_LOGIC);
END MINUTE;
ARCHITECTURE BEHAVE OF MINUTE IS
	SIGNAL COUNT1, COUNT0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN
	PROCESS (CLK)
	BEGIN
		IF (CLR = '0') THEN
			COUNT1 <= "0000";
			COUNT0 <= "0000";
		ELSIF (CLK'EVENT AND CLK = '1') THEN
			IF EN = '1' THEN
				IF COUNT1 = "0101" AND COUNT0 = "1001" THEN
					COUNT1 <= "0000";
					COUNT0 <= "0000";
					CO <= '1';
				ELSIF COUNT0 = "1001" THEN
					COUNT0 <= "0000";
					COUNT1 <= COUNT1 + '1';
				ELSE
					COUNT0 <= COUNT0 + '1';
					CO <= '0';
				END IF;
			END IF;
		END IF;
		MIN1 <= COUNT1;
		MIN0 <= COUNT0;
	END PROCESS;
END BEHAVE;