LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY DISPLAYDECOD IS
	PORT (
		NUM : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		DISPLAYOUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END DISPLAYDECOD;
ARCHITECTURE BEHAV OF DISPLAYDECOD IS
	SIGNAL DIS : STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN
	PROCESS (NUM)
	BEGIN
		CASE NUM IS
			WHEN "0000" => DIS <= "00111111";
			WHEN "0001" => DIS <= "00000110";
			WHEN "0010" => DIS <= "01011011";
			WHEN "0011" => DIS <= "01001111";
			WHEN "0100" => DIS <= "01100110";
			WHEN "0101" => DIS <= "01101101";
			WHEN "0110" => DIS <= "01111101";
			WHEN "0111" => DIS <= "00000111";
			WHEN "1000" => DIS <= "01111111";
			WHEN "1001" => DIS <= "01101111";
			WHEN "1111" => DIS <= "01000000";
			WHEN OTHERS => DIS <= "00000000";
		END CASE;
		DISPLAYOUT <= DIS;
	END PROCESS;
END BEHAV;