LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY DECODE138 IS
	PORT (
		DIN : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		DOUT : OUT STD_LOGIC_VECTOR (0 TO 7));
END DECODE138;
ARCHITECTURE BEHAV OF DECODE138 IS
BEGIN
	PROCESS (DIN)
	BEGIN
		IF (DIN = "111") THEN
			DOUT <= "11111110";
		ELSIF (DIN = "110") THEN
			DOUT <= "11111101";
		ELSIF (DIN = "101") THEN
			DOUT <= "11111011";
		ELSIF (DIN = "100") THEN
			DOUT <= "11110111";
		ELSIF (DIN = "011") THEN
			DOUT <= "11101111";
		ELSIF (DIN = "010") THEN
			DOUT <= "11011111";
		ELSIF (DIN = "001") THEN
			DOUT <= "10111111";
		ELSE
			DOUT <= "01111111";
		END IF;
	END PROCESS;
END BEHAV;